// AND Gate logic

module ANDGate (
	input wire A,B,
	output wire Cout);
	
	
	assign Cout = A & B;		// AND Gate operation
	
	endmodule
	
		

